* Testbench to show IV curves for an NMOS

*--------------------------------------------------------------
* INCLUDE
*--------------------------------------------------------------
.include ../../../lib/SUN_TRIO_GF130N.spi
.include ../../../models/ptm_130.spi

*--------------------------------------------------------------
* SOURCES
*--------------------------------------------------------------
vdrain D 0 dc 1
vgate G 0 dc 0.5

* Voltage source to make it easy to mesure current through transistor
vcur S 0 dc 0

*--------------------------------------------------------------
* DUT
*--------------------------------------------------------------
X1 D G S 0 NCHIO

*--------------------------------------------------------------
* ANALYSIS
*--------------------------------------------------------------
.dc vgate 0 1.8 0.1

*--------------------------------------------------------------
* CONTROL
*--------------------------------------------------------------
.control
run
plot ylog I(vcur)
.endc
.end
