* Equal strength

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../models/ptm_130.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20

.param p_vdd = 1.5
.param p_wp = 1
*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc p_vdd
V3 VSS 0 dc 0

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
M1 VG VG VSS VSS nmos W=0.65u L=0.13u
M2 VG VG VDD VDD pmos W={0.65u*p_wp} L=0.13u

*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
.op

.plot v(vg)
