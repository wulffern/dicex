
module mazeEscaper ( input [7:0][7:0] maze )

endmodule
