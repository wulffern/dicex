
module IVX1_CV(A, Y);
   input A;
   output Y;
endmodule // IVX1_CV

module BFX1_CV(A, Y);
   input A;
   output Y;
endmodule



module NDX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule


module ANX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule // ANX1_CV

module ORX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule // ORX1_CV

module EOX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule // EOX1_CV

module ENX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule





module NRX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule


module DFSRQNX1_CV(D,CK,S, R, Q, QN);
   input D,CK,S,R;
   output Q,QN;

endmodule
