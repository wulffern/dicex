* Check op

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20 reltol=1e-6 abstol=1e-8

.param sq={10}
.param l={0.15u}
.param w={sq*L}

.param In={60u}
.param Ip={In/6}


.param V_T = 25.9m
.param n = 1.5

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------

V2 VSS 0 dc 0
V1 VDD 0 dc 1.5
V3 VD 0 dc 1
V4 VG 0 dc 0.5

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------

*NMOS

M1 VD VG VSS VSS nmos W=w L=l

*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
*.dc I1 0.01u 10u 0.1u

.dc V4 0.4 0.6 0.01

*.dc I1  1p 1000u 100n

.defwave gmid_weak = 1/(n*V_T)
.defwave gmid_strong = 2/vgsteff(m1)
.defwave gmid = gm(m1)/id(m1)

.plot gm(m1) vt(m1) v(gmid_weak) v(gmid_strong) v(gmid) id(m1) vgsteff(m1)
