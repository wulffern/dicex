* Check op

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20 reltol=1e-6 abstol=1e-8

.param sq={10}
.param l={0.50u}
.param w={sq*L}

.param In={60u}
.param Ip={In/6}

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------

V2 VSS 0 dc 0
V1 VDD 0 dc 1.5

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------

*NMOS
I1 0 VDN dc In
M1 VDN VDN VSS VSS nmos W=w L=l

*PMOS
I2 VDP 0 dc Ip
M2 VDP VDP VDD VDD pmos W=w L=l

*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
.op
