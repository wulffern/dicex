
.SUBCKT NCHCM D G S B M=1 w=0.5u l=0.5u
M1 D G N1 B nmos W=w L=l
M2 N1  G N2 B nmos W=w L=l
M3 N2  G N3 B nmos W=w L=l
M4 N3  G N4 B nmos W=w L=l
M5 N4  G N5 B nmos W=w L=l
M6 N5  G S B nmos W=w L=l
.ends


.subckt CMIRR VDN IDN1 IDN2 IDN3 VSS

XM0 VDN VDN VSS VSS NCHCM

XM1a IDN1 VDN VSS VSS NCHCM
XM1b IDN1 VDN VSS VSS NCHCM

XM2a IDN2 VDN VSS VSS NCHCM
XM2b IDN2 VDN VSS VSS NCHCM
XM2c IDN2 VDN VSS VSS NCHCM
XM2d IDN2 VDN VSS VSS NCHCM

XM3a IDN3 VDN VSS VSS NCHCM
XM3b IDN3 VDN VSS VSS NCHCM
XM3c IDN3 VDN VSS VSS NCHCM
XM3d IDN3 VDN VSS VSS NCHCM
XM3e IDN3 VDN VSS VSS NCHCM
XM3f IDN3 VDN VSS VSS NCHCM
XM3g IDN3 VDN VSS VSS NCHCM
XM3h IDN3 VDN VSS VSS NCHCM


.ENDS
