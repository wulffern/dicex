module mazegen_tb;


   //------------------------------------------------------------
   // Testbench clock
   //------------------------------------------------------------
   logic clk =0;
   logic rst =0;
   int   cycles  =0 ;

   parameter integer clk_period = 1;
   parameter integer sim_end = clk_period*5000;
   always #clk_period clk=~clk;

   always @(posedge clk) begin
      if(cycles == 0)
        rst = 1;
      if(cycles == 1)
        rst = 0;
      cycles +=1;
   end


   logic [15:0] seed;
   parameter size = `MAZE_SIZE;
   parameter N = $clog2(size);

   tri [size-1:0] maze[size-1:0];
   tri             done;

   mazegen #(.size(size),.N(N)) mz(clk,rst,seed,done,maze);

   //------------------------------------------------------------
   // Testbench stuff
   //------------------------------------------------------------
   int                   fd,fo,fp;
   int                   idx;
   int                   str;
   int                x,y;

   initial
     begin

        seed = `MAZE_SEED;

        $dumpfile("mazegen_tb.vcd");
        $dumpvars(0,mazegen_tb);


        fo = $fopen("maze.txt","w");
        #sim_end
          for (y = 0; y<size; y=y+1) begin
               $fwrite(fo,"%b\n",maze[y]);
          end

        #sim_end $fclose(fo);

        #sim_end
          $stop;



     end

endmodule
