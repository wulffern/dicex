
module mazeEscaper ( input [7:0] maze [7:0],
                     input        startX [7:0],
                     input        startY [7:0],
                     input        clk,
                     input        reset,
                     output [7:0] path [7:0]);

endmodule
