* Check op

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20 reltol=1e-6 abstol=1e-8

.param sq={10}
.param l={0.50u}
.param w={sq*L}

.param In={10u}
.param Ip={In/6}

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------

V2 VSS 0 dc 0
V1 VDD 0 dc 1.5

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------

*NMOS
I1 0 VDN dc In
M1 VDN VDN N1 VSS nmos W=w L=l
M2 N1  VDN N2 VSS nmos W=w L=l
M3 N2  VDN N3 VSS nmos W=w L=l
M4 N3  VDN N4 VSS nmos W=w L=l
M5 N4  VDN N5 VSS nmos W=w L=l
M6 N5  VDN VSS VSS nmos W=w L=l


*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
.op
