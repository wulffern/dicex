* Gate Voltage sweep

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../models/ptm_130.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
V1 VD VSS dc 1.5
V2 VG VSS dc 0
V3 VSS 0 dc 0

.param k_weak=0.04m
.param k_strong=3.9m
.param k_sat=1.5m
.param n = 1.5
.param V_T = 25.6m


*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
M1 VD VG VSS VSS nmos W=2u L=0.2u

*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
.dc V2 0 1.5 0.01
.defwave a = gm(m1)*rds(m1)
.defwave id_weak = k_weak*exp(vgt(m1)/(n*V_T))
.defwave id_strong = k_strong*vgsteff(m1)*vgsteff(m1) + k_weak
.defwave id_sat = k_sat*vgt(m1)

.plot v(vg) gm(m1) rds(m1) id(m1) v(a) q(id_weak) v(id_strong) v(id_sat)
