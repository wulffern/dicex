.SUBCKT PCHIO D G S B
M1 D G S B pmos  w=1.08u  l=0.6u
.ENDS

.SUBCKT NCHIO D G S B
M1 D G S B nmos  w=1.08u  l=0.6u
.ENDS

.SUBCKT NCHIOCM D G S B
XM0 N0 G S B NCHIO 
XM1 N1 G N0 B NCHIO 
XM4 N2 G N1 B NCHIO 
XM5 D G N2 B NCHIO 
.ENDS

.SUBCKT PCHIOCM D G S B
XM0 N0 G S B PCHIO 
XM1 N1 G N0 B PCHIO 
XM4 N2 G N1 B PCHIO 
XM5 D G N2 B PCHIO 
.ENDS

.SUBCKT NCHIOA D G S B
XM0 D G S B NCHIO 
XM1 S G D B NCHIO 
.ENDS

.SUBCKT PCHIOA D G S B
XM0 D G S B PCHIO 
XM1 S G D B PCHIO 
.ENDS

.SUBCKT NCHIOCM2 D G S B
XM0 D G S B NCHIOCM 
XM1 S G D B NCHIOCM 
.ENDS

.SUBCKT PCHIOCM2 D G S B
XM0 D G S B PCHIOCM 
XM1 S G D B PCHIOCM 
.ENDS

.SUBCKT PCHIO_4C D G S B
M1 D G S B pmos  w=2.52u  l=0.6u
.ENDS

.SUBCKT PCHIOA_4C D G S B
XM0 D G S B PCHIO_4C 
XM1 S G D B PCHIO_4C 
.ENDS

.SUBCKT PCHIOCM_4C D G S B
XM0 N0 G S B PCHIO_4C 
XM1 N1 G N0 B PCHIO_4C 
XM4 N2 G N1 B PCHIO_4C 
XM5 D G N2 B PCHIO_4C 
.ENDS

.SUBCKT PCHIOCM2_4C D G S B
XM0 D G S B PCHIOCM_4C 
XM1 S G D B PCHIOCM_4C 
.ENDS

.SUBCKT PCHIO_6C D G S B
M1 D G S B pmos  w=3.96u  l=0.6u
.ENDS

.SUBCKT PCHIOA_6C D G S B
XM0 D G S B PCHIO_6C 
XM1 S G D B PCHIO_6C 
.ENDS

.SUBCKT PCHIOCM_6C D G S B
XM0 N0 G S B PCHIO_6C 
XM1 N1 G N0 B PCHIO_6C 
XM4 N2 G N1 B PCHIO_6C 
XM5 D G N2 B PCHIO_6C 
.ENDS

.SUBCKT PCHIOCM2_6C D G S B
XM0 D G S B PCHIOCM_6C 
XM1 S G D B PCHIOCM_6C 
.ENDS

.SUBCKT PCHIO_10C D G S B
M1 D G S B pmos  w=6.84u  l=0.6u
.ENDS

.SUBCKT PCHIOA_10C D G S B
XM0 D G S B PCHIO_10C 
XM1 S G D B PCHIO_10C 
.ENDS

.SUBCKT PCHIOCM_10C D G S B
XM0 N0 G S B PCHIO_10C 
XM1 N1 G N0 B PCHIO_10C 
XM4 N2 G N1 B PCHIO_10C 
XM5 D G N2 B PCHIO_10C 
.ENDS

.SUBCKT PCHIOCM2_10C D G S B
XM0 D G S B PCHIOCM_10C 
XM1 S G D B PCHIOCM_10C 
.ENDS

.SUBCKT PCHIO_12C D G S B
M1 D G S B pmos  w=8.28u  l=0.6u
.ENDS

.SUBCKT PCHIOA_12C D G S B
XM0 D G S B PCHIO_12C 
XM1 S G D B PCHIO_12C 
.ENDS

.SUBCKT PCHIOCM_12C D G S B
XM0 N0 G S B PCHIO_12C 
XM1 N1 G N0 B PCHIO_12C 
XM4 N2 G N1 B PCHIO_12C 
XM5 D G N2 B PCHIO_12C 
.ENDS

.SUBCKT PCHIOCM2_12C D G S B
XM0 D G S B PCHIOCM_12C 
XM1 S G D B PCHIOCM_12C 
.ENDS

.SUBCKT NCHIO_4C D G S B
M1 D G S B nmos  w=2.52u  l=0.6u
.ENDS

.SUBCKT NCHIOA_4C D G S B
XM0 D G S B NCHIO_4C 
XM1 S G D B NCHIO_4C 
.ENDS

.SUBCKT NCHIOCM_4C D G S B
XM0 N0 G S B NCHIO_4C 
XM1 N1 G N0 B NCHIO_4C 
XM4 N2 G N1 B NCHIO_4C 
XM5 D G N2 B NCHIO_4C 
.ENDS

.SUBCKT NCHIOCM2_4C D G S B
XM0 D G S B NCHIOCM_4C 
XM1 S G D B NCHIOCM_4C 
.ENDS

.SUBCKT NCHIO_6C D G S B
M1 D G S B nmos  w=3.96u  l=0.6u
.ENDS

.SUBCKT NCHIOA_6C D G S B
XM0 D G S B NCHIO_6C 
XM1 S G D B NCHIO_6C 
.ENDS

.SUBCKT NCHIOCM_6C D G S B
XM0 N0 G S B NCHIO_6C 
XM1 N1 G N0 B NCHIO_6C 
XM4 N2 G N1 B NCHIO_6C 
XM5 D G N2 B NCHIO_6C 
.ENDS

.SUBCKT NCHIOCM2_6C D G S B
XM0 D G S B NCHIOCM_6C 
XM1 S G D B NCHIOCM_6C 
.ENDS

.SUBCKT NCHIO_10C D G S B
M1 D G S B nmos  w=6.84u  l=0.6u
.ENDS

.SUBCKT NCHIOA_10C D G S B
XM0 D G S B NCHIO_10C 
XM1 S G D B NCHIO_10C 
.ENDS

.SUBCKT NCHIOCM_10C D G S B
XM0 N0 G S B NCHIO_10C 
XM1 N1 G N0 B NCHIO_10C 
XM4 N2 G N1 B NCHIO_10C 
XM5 D G N2 B NCHIO_10C 
.ENDS

.SUBCKT NCHIOCM2_10C D G S B
XM0 D G S B NCHIOCM_10C 
XM1 S G D B NCHIOCM_10C 
.ENDS

.SUBCKT NCHIO_12C D G S B
M1 D G S B nmos  w=8.28u  l=0.6u
.ENDS

.SUBCKT NCHIOA_12C D G S B
XM0 D G S B NCHIO_12C 
XM1 S G D B NCHIO_12C 
.ENDS

.SUBCKT NCHIOCM_12C D G S B
XM0 N0 G S B NCHIO_12C 
XM1 N1 G N0 B NCHIO_12C 
XM4 N2 G N1 B NCHIO_12C 
XM5 D G N2 B NCHIO_12C 
.ENDS

.SUBCKT NCHIOCM2_12C D G S B
XM0 D G S B NCHIOCM_12C 
XM1 S G D B NCHIOCM_12C 
.ENDS

.SUBCKT TAPCELLB_EV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS NCHIO 
XMP1 AVDD AVDD AVDD AVDD PCHIO 
.ENDS

.SUBCKT TIEH_EV Y AVDD AVSS
XMN0 A A AVSS AVSS NCHIO 
XMP0 Y A AVDD AVDD PCHIO 
.ENDS

.SUBCKT TIEL_EV Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMP0 A A AVDD AVDD PCHIO 
.ENDS

.SUBCKT IVX1_EV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMP0 Y A AVDD AVDD PCHIO 
.ENDS

.SUBCKT IVX2_EV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMN1 AVSS A Y AVSS NCHIO 
XMP0 Y A AVDD AVDD PCHIO 
XMP1 AVDD A Y AVDD PCHIO 
.ENDS

.SUBCKT IVX4_EV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMN1 AVSS A Y AVSS NCHIO 
XMN2 Y A AVSS AVSS NCHIO 
XMN3 AVSS A Y AVSS NCHIO 
XMP0 Y A AVDD AVDD PCHIO 
XMP1 AVDD A Y AVDD PCHIO 
XMP2 Y A AVDD AVDD PCHIO 
XMP3 AVDD A Y AVDD PCHIO 
.ENDS

.SUBCKT IVX8_EV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMN1 AVSS A Y AVSS NCHIO 
XMN2 Y A AVSS AVSS NCHIO 
XMN3 AVSS A Y AVSS NCHIO 
XMN4 Y A AVSS AVSS NCHIO 
XMN5 AVSS A Y AVSS NCHIO 
XMN6 Y A AVSS AVSS NCHIO 
XMN7 AVSS A Y AVSS NCHIO 
XMP0 Y A AVDD AVDD PCHIO 
XMP1 AVDD A Y AVDD PCHIO 
XMP2 Y A AVDD AVDD PCHIO 
XMP3 AVDD A Y AVDD PCHIO 
XMP4 Y A AVDD AVDD PCHIO 
XMP5 AVDD A Y AVDD PCHIO 
XMP6 Y A AVDD AVDD PCHIO 
XMP7 AVDD A Y AVDD PCHIO 
.ENDS

.SUBCKT BFX1_EV A Y AVDD AVSS
XMN0 AVSS A B AVSS NCHIO 
XMN1 Y B AVSS AVSS NCHIO 
XMP0 AVDD A B AVDD PCHIO 
XMP1 Y B AVDD AVDD PCHIO 
.ENDS

.SUBCKT NRX1_EV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMN1 AVSS B Y AVSS NCHIO 
XMP0 N1 A AVDD AVDD PCHIO 
XMP1 Y B N1 AVDD PCHIO 
.ENDS

.SUBCKT NDX1_EV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS NCHIO 
XMN1 Y B N1 AVSS NCHIO 
XMP0 Y A AVDD AVDD PCHIO 
XMP1 AVDD B Y AVDD PCHIO 
.ENDS

.SUBCKT ORX1_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT ORX2_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT ORX4_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT ANX1_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT ANX2_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT ANX4_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT ANX8_EV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_EV 
XA2 YN Y AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT IVTRIX1_EV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS NCHIO 
XMN1 Y C N1 AVSS NCHIO 
XMP0 N2 A AVDD AVDD PCHIO 
XMP1 Y CN N2 AVDD PCHIO 
.ENDS

.SUBCKT NDTRIX1_EV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS NCHIO 
XMN0 N2 A N1 AVSS NCHIO 
XMN1 Y C N2 AVSS NCHIO 
XMP2 AVDD RN N2 AVDD PCHIO 
XMP0 N2 A AVDD AVDD PCHIO 
XMP1 Y CN N2 AVDD PCHIO 
.ENDS

.SUBCKT DFRNQNX1_EV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_EV 
XA1 CK RN CKN AVDD AVSS NDX1_EV 
XA2 CKN CKB AVDD AVSS IVX1_EV 
XA3 D CKN CKB A0 AVDD AVSS IVTRIX1_EV 
XA4 A1 CKB CKN A0 AVDD AVSS IVTRIX1_EV 
XA5 A0 A1 AVDD AVSS IVX1_EV 
XA6 A1 CKB CKN QN AVDD AVSS IVTRIX1_EV 
XA7 Q CKN CKB RN QN AVDD AVSS NDTRIX1_EV 
XA8 QN Q AVDD AVSS IVX1_EV 
.ENDS

.SUBCKT SCX1_EV A Y AVDD AVSS
XA2 N1 A AVSS AVSS NCHIO 
XA3 SCO A N1 AVSS NCHIO 
XA4a AVDD SCO N1 AVSS NCHIO 
XA4b AVDD SCO N1 AVSS NCHIO 
XA5 Y SCO AVSS AVSS NCHIO 
XB0 N2 A AVDD AVDD PCHIO 
XB1 SCO A N2 AVDD PCHIO 
XB3a N2 SCO AVSS AVDD PCHIO 
XB3b N2 SCO AVSS AVDD PCHIO 
XB4 Y SCO AVDD AVDD PCHIO 
.ENDS

.SUBCKT SWX2_EV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMN1 AVSS A Y AVSS NCHIO 
XMP0 Y A VREF AVDD PCHIO 
XMP1 VREF A Y AVDD PCHIO 
.ENDS

.SUBCKT SWX4_EV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS NCHIO 
XMN1 AVSS A Y AVSS NCHIO 
XMN2 Y A AVSS AVSS NCHIO 
XMN3 AVSS A Y AVSS NCHIO 
XMP0 Y A VREF AVDD PCHIO 
XMP1 VREF A Y AVDD PCHIO 
XMP2 Y A VREF AVDD PCHIO 
XMP3 VREF A Y AVDD PCHIO 
.ENDS

.SUBCKT TGPD_EV C A B AVDD AVSS
XMN0 AVSS C CN AVSS NCHIO 
XMN1 B C AVSS AVSS NCHIO 
XMN2 A CN B AVSS NCHIO 
XMP0 AVDD C CN AVDD PCHIO 
XMP1_DMY B AVDD AVDD AVDD PCHIO 
XMP2 A C B AVDD PCHIO 
.ENDS

.SUBCKT SUN_TRIO AVDD AVSS
XA0 AVDD AVSS TAPCELLB_EV 
XA1 Y1 AVDD AVSS TIEH_EV 
XA2 Y2 AVDD AVSS TIEL_EV 
XB0 AVDD AVSS TAPCELLB_EV 
XB3 A3 Y3 AVDD AVSS IVX1_EV 
XB4 A4 Y4 AVDD AVSS IVX2_EV 
XB5 A5 Y5 AVDD AVSS IVX4_EV 
XB6 A6 Y6 AVDD AVSS IVX8_EV 
XC0 AVDD AVSS TAPCELLB_EV 
XC7 A7 Y7 AVDD AVSS BFX1_EV 
XD0 AVDD AVSS TAPCELLB_EV 
XD8 A8 B8 Y8 AVDD AVSS NRX1_EV 
XD9 A9 B9 Y9 AVDD AVSS NDX1_EV 
XD10 A10 B10 Y10 AVDD AVSS ORX1_EV 
XD11 A11 B11 Y11 AVDD AVSS ANX1_EV 
XE0 AVDD AVSS TAPCELLB_EV 
XE12 A12 Y12 AVDD AVSS SCX1_EV 
XF0 AVDD AVSS TAPCELLB_EV 
XF13 A13 Y13 V13 AVDD AVSS SWX2_EV 
XF14 A14 Y14 V14 AVDD AVSS SWX4_EV 
XF15 A15 Y15 V15 AVDD AVSS TGPD_EV 
.ENDS

