* Check op

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20 reltol=1e-6 abstol=1e-8

.param sq={10}
.param l={0.15u}
.param w={sq*L}

.param In={60u}
.param Ip={In/6}


.param V_T = 25.9m
.param n = 1.5

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------

V2 VSS 0 dc 0
V1 VDD 0 dc 1.5

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------

*NMOS
I1 0 VDN dc In
M1 VDN VDN VSS VSS nmos W=w L=l

*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
*.dc I1 0.01u 2u 0.1u

.dc I1 50u 1000u 0.1u

*.dc I1  1p 1000u 100n

.defwave gmid_weak = 1/(n*V_T)
.defwave gmid_strong = 2/vgt(m1)
.defwave gmid = gm(m1)/id(m1)

.plot gm(m1) vt(m1) v(gmid_weak) v(gmid_strong) v(gmid)
