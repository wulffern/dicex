
module IVX1_CV(A, Y);
   input A;
   output Y;
endmodule


module NDX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule


module NRX1_CV(A, B, Y);
   input A,B;
   output Y;
endmodule


module DFSRQNX1_CV(D,CK,S, R, Q, QN);
   input D,CK,S,R;
   output Q,QN;

endmodule
