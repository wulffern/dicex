
.SUBCKT PIXEL_SENSOR VBN1 VBN2 RAMP RESET ERASE EXPOSE READ
+ DATA[7] DATA[6] DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0]

.ENDS
