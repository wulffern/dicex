
.subckt OTA VIP VIN VO VDD VSS IBP

MP1 VDP VDP VDD VDD pmos L=0.5u W=0.5u
MP2 VO VDP VDD VDD pmos L=0.5u W=0.5u

MN1 VO VIN VS VSS nmos L=0.15u W=0.5u
MN2 VDP VIP VS VSS nmos L=0.15u W=0.5u

XMN3 VS IBP VSS VSS NCHCM
XMN4 IBP IBP VSS VSS NCHCM

.ends
