* Transistor library

.SUBCKT PCH D G S B
M1 D G S B pmos  w=1.08u  l=0.13u
.ENDS

.SUBCKT NCH D G S B
M1 D G S B nmos  w=1.08u  l=0.13u
.ENDS

.SUBCKT NCHCM D G S B
XM0 N0 G S B NCH
XM1 N1 G N0 B NCH
XM4 N2 G N1 B NCH
XM5 D G N2 B NCH
.ENDS

.SUBCKT PCHCM D G S B
XM0 N0 G S B PCH
XM1 N1 G N0 B PCH
XM4 N2 G N1 B PCH
XM5 D G N2 B PCH
.ENDS

.SUBCKT NCHA D G S B
XM0 D G S B NCH
XM1 S G D B NCH
.ENDS

.SUBCKT PCHA D G S B
XM0 D G S B PCH
XM1 S G D B PCH
.ENDS

.SUBCKT NCHCM2 D G S B
XM0 D G S B NCHCM
XM1 S G D B NCHCM
.ENDS

.SUBCKT PCHCM2 D G S B
XM0 D G S B PCHCM
XM1 S G D B PCHCM
.ENDS

.SUBCKT PCH_4C D G S B
M1 D G S B pmos  w=2.52u  l=0.13u
.ENDS

.SUBCKT PCHA_4C D G S B
XM0 D G S B PCH_4C
XM1 S G D B PCH_4C
.ENDS

.SUBCKT PCHCM_4C D G S B
XM0 N0 G S B PCH_4C
XM1 N1 G N0 B PCH_4C
XM4 N2 G N1 B PCH_4C
XM5 D G N2 B PCH_4C
.ENDS

.SUBCKT PCHCM2_4C D G S B
XM0 D G S B PCHCM_4C
XM1 S G D B PCHCM_4C
.ENDS

.SUBCKT PCH_6C D G S B
M1 D G S B pmos  w=3.96u  l=0.13u
.ENDS

.SUBCKT PCHA_6C D G S B
XM0 D G S B PCH_6C
XM1 S G D B PCH_6C
.ENDS

.SUBCKT PCHCM_6C D G S B
XM0 N0 G S B PCH_6C
XM1 N1 G N0 B PCH_6C
XM4 N2 G N1 B PCH_6C
XM5 D G N2 B PCH_6C
.ENDS

.SUBCKT PCHCM2_6C D G S B
XM0 D G S B PCHCM_6C
XM1 S G D B PCHCM_6C
.ENDS

.SUBCKT PCH_10C D G S B
M1 D G S B pmos  w=6.84u  l=0.13u
.ENDS

.SUBCKT PCHA_10C D G S B
XM0 D G S B PCH_10C
XM1 S G D B PCH_10C
.ENDS

.SUBCKT PCHCM_10C D G S B
XM0 N0 G S B PCH_10C
XM1 N1 G N0 B PCH_10C
XM4 N2 G N1 B PCH_10C
XM5 D G N2 B PCH_10C
.ENDS

.SUBCKT PCHCM2_10C D G S B
XM0 D G S B PCHCM_10C
XM1 S G D B PCHCM_10C
.ENDS

.SUBCKT PCH_12C D G S B
M1 D G S B pmos  w=8.28u  l=0.13u
.ENDS

.SUBCKT PCHA_12C D G S B
XM0 D G S B PCH_12C
XM1 S G D B PCH_12C
.ENDS

.SUBCKT PCHCM_12C D G S B
XM0 N0 G S B PCH_12C
XM1 N1 G N0 B PCH_12C
XM4 N2 G N1 B PCH_12C
XM5 D G N2 B PCH_12C
.ENDS

.SUBCKT PCHCM2_12C D G S B
XM0 D G S B PCHCM_12C
XM1 S G D B PCHCM_12C
.ENDS

.SUBCKT NCH_4C D G S B
M1 D G S B nmos  w=2.52u  l=0.13u
.ENDS

.SUBCKT NCHA_4C D G S B
XM0 D G S B NCH_4C
XM1 S G D B NCH_4C
.ENDS

.SUBCKT NCHCM_4C D G S B
XM0 N0 G S B NCH_4C
XM1 N1 G N0 B NCH_4C
XM4 N2 G N1 B NCH_4C
XM5 D G N2 B NCH_4C
.ENDS

.SUBCKT NCHCM2_4C D G S B
XM0 D G S B NCHCM_4C
XM1 S G D B NCHCM_4C
.ENDS

.SUBCKT NCH_6C D G S B
M1 D G S B nmos  w=3.96u  l=0.13u
.ENDS

.SUBCKT NCHA_6C D G S B
XM0 D G S B NCH_6C
XM1 S G D B NCH_6C
.ENDS

.SUBCKT NCHCM_6C D G S B
XM0 N0 G S B NCH_6C
XM1 N1 G N0 B NCH_6C
XM4 N2 G N1 B NCH_6C
XM5 D G N2 B NCH_6C
.ENDS

.SUBCKT NCHCM2_6C D G S B
XM0 D G S B NCHCM_6C
XM1 S G D B NCHCM_6C
.ENDS

.SUBCKT NCH_10C D G S B
M1 D G S B nmos  w=6.84u  l=0.13u
.ENDS

.SUBCKT NCHA_10C D G S B
XM0 D G S B NCH_10C
XM1 S G D B NCH_10C
.ENDS

.SUBCKT NCHCM_10C D G S B
XM0 N0 G S B NCH_10C
XM1 N1 G N0 B NCH_10C
XM4 N2 G N1 B NCH_10C
XM5 D G N2 B NCH_10C
.ENDS

.SUBCKT NCHCM2_10C D G S B
XM0 D G S B NCHCM_10C
XM1 S G D B NCHCM_10C
.ENDS

.SUBCKT NCH_12C D G S B
M1 D G S B nmos  w=8.28u  l=0.13u
.ENDS

.SUBCKT NCHA_12C D G S B
XM0 D G S B NCH_12C
XM1 S G D B NCH_12C
.ENDS

.SUBCKT NCHCM_12C D G S B
XM0 N0 G S B NCH_12C
XM1 N1 G N0 B NCH_12C
XM4 N2 G N1 B NCH_12C
XM5 D G N2 B NCH_12C
.ENDS

.SUBCKT NCHCM2_12C D G S B
XM0 D G S B NCHCM_12C
XM1 S G D B NCHCM_12C
.ENDS

.SUBCKT TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS NCH
XMP1 AVDD AVDD AVDD AVDD PCH
.ENDS

.SUBCKT TIEH_CV Y AVDD AVSS
XMN0 A A AVSS AVSS NCH
XMP0 Y A AVDD AVDD PCH
.ENDS

.SUBCKT TIEL_CV Y AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMP0 A A AVDD AVDD PCH
.ENDS

.SUBCKT IVX1_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMP0 Y A AVDD AVDD PCH
.ENDS

.SUBCKT IVX2_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMN1 AVSS A Y AVSS NCH
XMP0 Y A AVDD AVDD PCH
XMP1 AVDD A Y AVDD PCH
.ENDS

.SUBCKT IVX4_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMN1 AVSS A Y AVSS NCH
XMN2 Y A AVSS AVSS NCH
XMN3 AVSS A Y AVSS NCH
XMP0 Y A AVDD AVDD PCH
XMP1 AVDD A Y AVDD PCH
XMP2 Y A AVDD AVDD PCH
XMP3 AVDD A Y AVDD PCH
.ENDS

.SUBCKT IVX8_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMN1 AVSS A Y AVSS NCH
XMN2 Y A AVSS AVSS NCH
XMN3 AVSS A Y AVSS NCH
XMN4 Y A AVSS AVSS NCH
XMN5 AVSS A Y AVSS NCH
XMN6 Y A AVSS AVSS NCH
XMN7 AVSS A Y AVSS NCH
XMP0 Y A AVDD AVDD PCH
XMP1 AVDD A Y AVDD PCH
XMP2 Y A AVDD AVDD PCH
XMP3 AVDD A Y AVDD PCH
XMP4 Y A AVDD AVDD PCH
XMP5 AVDD A Y AVDD PCH
XMP6 Y A AVDD AVDD PCH
XMP7 AVDD A Y AVDD PCH
.ENDS

.SUBCKT BFX1_CV A Y AVDD AVSS
XMN0 AVSS A B AVSS NCH
XMN1 Y B AVSS AVSS NCH
XMP0 AVDD A B AVDD PCH
XMP1 Y B AVDD AVDD PCH
.ENDS

.SUBCKT NRX1_CV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMN1 AVSS B Y AVSS NCH
XMP0 N1 A AVDD AVDD PCH
XMP1 Y B N1 AVDD PCH
.ENDS

.SUBCKT NDX1_CV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS NCH
XMN1 Y B N1 AVSS NCH
XMP0 Y A AVDD AVDD PCH
XMP1 AVDD B Y AVDD PCH
.ENDS

.SUBCKT ORX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ORX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ORX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX8_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT IVTRIX1_CV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS NCH
XMN1 Y C N1 AVSS NCH
XMP0 N2 A AVDD AVDD PCH
XMP1 Y CN N2 AVDD PCH
.ENDS

.SUBCKT NDTRIX1_CV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS NCH
XMN0 N2 A N1 AVSS NCH
XMN1 Y C N2 AVSS NCH
XMP2 AVDD RN N2 AVDD PCH
XMP0 N2 A AVDD AVDD PCH
XMP1 Y CN N2 AVDD PCH
.ENDS

.SUBCKT DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS IVTRIX1_CV
XA5 A0 A1 AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS NDTRIX1_CV
XA8 QN Q AVDD AVSS IVX1_CV
.ENDS


.SUBCKT DFSRQNX1_CV D CK S R Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA0a R RN AVDD AVSS IVX1_CV
XA1 CK RN CKN AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS IVTRIX1_CV
XA5 A0 A1 AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS NDTRIX1_CV
XA8 QN Q AVDD AVSS IVX1_CV
.ENDS



.SUBCKT SCX1_CV A Y AVDD AVSS
XA2 N1 A AVSS AVSS NCH
XA3 SCO A N1 AVSS NCH
XA4a AVDD SCO N1 AVSS NCH
XA4b AVDD SCO N1 AVSS NCH
XA5 Y SCO AVSS AVSS NCH
XB0 N2 A AVDD AVDD PCH
XB1 SCO A N2 AVDD PCH
XB3a N2 SCO AVSS AVDD PCH
XB3b N2 SCO AVSS AVDD PCH
XB4 Y SCO AVDD AVDD PCH
.ENDS

.SUBCKT SWX2_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMN1 AVSS A Y AVSS NCH
XMP0 Y A VREF AVDD PCH
XMP1 VREF A Y AVDD PCH
.ENDS

.SUBCKT SWX4_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS NCH
XMN1 AVSS A Y AVSS NCH
XMN2 Y A AVSS AVSS NCH
XMN3 AVSS A Y AVSS NCH
XMP0 Y A VREF AVDD PCH
XMP1 VREF A Y AVDD PCH
XMP2 Y A VREF AVDD PCH
XMP3 VREF A Y AVDD PCH
.ENDS

.SUBCKT TGPD_CV C A B AVDD AVSS
XMN0 AVSS C CN AVSS NCH
XMN1 B C AVSS AVSS NCH
XMN2 A CN B AVSS NCH
XMP0 AVDD C CN AVDD PCH
XMP1_DMY B AVDD AVDD AVDD PCH
XMP2 A C B AVDD PCH
.ENDS

.SUBCKT SUN_TR AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 Y1 AVDD AVSS TIEH_CV
XA2 Y2 AVDD AVSS TIEL_CV
XB0 AVDD AVSS TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS IVX1_CV
XB4 A4 Y4 AVDD AVSS IVX2_CV
XB5 A5 Y5 AVDD AVSS IVX4_CV
XB6 A6 Y6 AVDD AVSS IVX8_CV
XC0 AVDD AVSS TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS BFX1_CV
XD0 AVDD AVSS TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS ANX1_CV
XE0 AVDD AVSS TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SCX1_CV
XF0 AVDD AVSS TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS TGPD_CV
.ENDS

